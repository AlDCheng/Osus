library verilog;
use verilog.vl_types.all;
entity image_process_tf is
end image_process_tf;

module test_rom(input wire [17:0] addr,
               input wire clk,
               output reg dout);
   // let the tools infer the right number of BRAMs
   //(* ram_style = "block" *)
   wire [587:0] mem;
   assign mem = 588'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111000000000000000000001111111100000000000000000001111111111000000000000000000111111111100000000000000000011111111110000000000000000001111111111000000000000000000011111111000000000000000000001111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
   
   always @(posedge clk) begin
     // if (we) mem[addr] <= din;
     if (addr < 588) dout <= mem[addr];
     else dout <= 0;
   end
endmodule
module mybram (input wire [9:0] addr,
               input wire clk,
               input wire din,
               output reg dout,
               input wire we);
   wire [615:0] mem;
   assign mem = 616'b0000000000000000000000010000001000000000000000000000000001000000000000000100000000001100000000000100011000000100100000001000000001000000010010000000000000000000000000001000100000000000000110000000100000000000001000111100000010000000001000000011010000001000000000000000000110000000100000000000000000000000000010000001100000000000000000000000001111100000000000000000000001111111000000011000100000000111111100000000000000000000011111110000000000000000000000111110000001000000100000100001110000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000;
   
   always @(posedge clk) begin
     // if (we) mem[addr] <= din;
     dout <= mem[addr];
   end
endmodule
